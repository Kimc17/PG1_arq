module TOP(input logic clk, reset);
logic [31:0] Inst, pc4, BranchDir, PC4, INST, ImmExtend, Data1, Data2,
DATA1, DATA2, IMMEXTEND, ALUResult, ALURESULT, DATA21, DATA5, ALURESULT2, DATA52, DataInput,
Data52;

logic WE,DataInputS, OpbSelect, RWrite, RWRITE, RWRITE2, RWRITE3, Branch, PCSelect,DataInputON,
 DATAINPUTON1, WE1, DATAINPUTS1, OPBSELECT, SELECTMEM1, SelectMem, 
 DATAINPUTON2,WE2, DATAINPUTS2, SELECTMEM2, DATAINPUTS3, DATAINPUTON3;
 
logic [2:0] ALUSignal, ALUSIGNAL ; 
logic [3:0] RD;

FETCH fetch(PCSelect, clk, reset, pc4, BranchDir, Inst, PC4);

REGFETCH rfetch(Inst, PC4, clk, reset, INST, pc4);


UNIDAD_CONTROL controlp( INST[31:27], INST[14:12], WE,DataInputS,
 DataInputON, OpbSelect, RWrite, Branch, SelectMem, ALUSignal);

DECO deco(INST[22:19], INST[18:15], INST[26:23],Branch, clk, DATAINPUTON3, RWrite, INST[18:0], DataInput, 
PCSelect, BranchDir, ImmExtend, Data1, Data2, RD );	 
 
REGDECO rdeco(Data1, Data2, ImmExtend,  DataInputON,clk, reset, WE, DataInputS, ALUSignal, OpbSelect, SelectMem,
DATAINPUTON1, DATA1, DATA2, IMMEXTEND, WE1, DATAINPUTS1, ALUSIGNAL, OPBSELECT, SELECTMEM1 );					 


EXE exe(IMMEXTEND, DATA2, DATA1, ALUSIGNAL, OPBSELECT, ALUResult);

REGEXE rexe(ALUResult, DATA2, DATAINPUTON1,clk, reset, WE1, DATAINPUTS1, SELECTMEM1,
ALURESULT, DATA21, DATAINPUTON2,WE2, DATAINPUTS2, SELECTMEM2 );

MEM mem(SELECTMEM2 , WE2, clk, ALURESULT, DATA21, DATA5);

REGMEM rmem(ALURESULT, DATA5, clk, reset, DATAINPUTON2, DATAINPUTS2, ALURESULT2, DATA52,DATAINPUTS3, DATAINPUTON3);

WB wbp(DATAINPUTS3, DATA52, ALURESULT2, DataInput);

endmodule